library verilog;
use verilog.vl_types.all;
entity Interpolador_vlg_vec_tst is
end Interpolador_vlg_vec_tst;
