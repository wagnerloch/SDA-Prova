library verilog;
use verilog.vl_types.all;
entity Upsampling_vlg_vec_tst is
end Upsampling_vlg_vec_tst;
